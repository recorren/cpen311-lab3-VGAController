library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.NbitRegDecs.all;

--Screen clearer module, runs an internal state machine on the rising edge of rst
--done is set to 1 after screen clear is complete. 

entity scrn_clearer is
  port(CLOCK_50: in std_logic;
       rst : in std_logic;
       color: out std_logic_vector(2 downto 0);
       x : out std_logic_vector(7 downto 0);
       y : out std_logic_vector(6 downto 0);
       plot : out std_logic;
       done : out std_logic);
end entity; 

architecture impl of scrn_clearer is
  
  signal currentX, nextX : std_logic_vector(x'LENGTH downto 0) := (others => '0'); 
  signal currentY, nextY : std_logic_vector(y'LENGTH downto 0) := (others => '0'); 
  signal xEqualsLimit : std_logic := '0'; 
  signal yEqualsLimit : std_logic := '0'; 

  begin
    --XPOS asynchronously resets to value 0 if rst is high
    
    XPOS : NbitReg generic map(x'LENGTH, 0)
                   port map(D => nextX, clk => CLOCK_50, Q => currentX, rst => rst);
    
    YPOS : NbitReg generic map(y'LENGTH, 0)
                   port map(D => nextY, clk => CLOCK_50, Q => currentY, rst => rst);
                     
    process(all) begin
      
    end process; 
    
end impl;